* AD8220 SPICE Macro-model               09/09, Rev. C
*                                        PRB IAP ADI
*
* Revision History:
* 
* Node assignments
*                 inverting input
*                 |   RG
*                 |   |    RG
*                 |   |    |  non_inverting input
*                 |   |    |    |    negative supply
*                 |   |    |    |    |    ref
*                 |   |    |    |    |    |   output
*                 |   |    |    |    |    |    |     positive supply
*                 |   |    |    |    |    |    |     |
.SUBCKT AD8220  IN-  RG-  RG+  IN+  -Vs   REF  VOUT  +Vs          
** INPUT STAGE
R1 N009 N008 20E3
R2 N008 Inverting_Out 20E3
R3 N013 noninverting_out 20.002e3
R4 REF N013 20e3
R5 RG- N003 24700
R6 RG+ N012 24724
D3 N003 P001 D
D4 P002 N003 D
V3 P002 VNEGx 0.84
V4 VPOSx P001 2.35
D5 N012 P003 D
D6 P004 N012 D
V5 P004 VNEGx 0.84
V6 VPOSx P003 2.35
D7 N005 P005 D
D8 P006 N005 D
V7 P006 VNEGx -10
V8 VPOSx P005 -10
D9 N019 P007 D
D10 P008 N019 D
V9 P008 VNEGx -10
V10 VPOSx P007 -10
D11 N009 P009 D
D12 P010 N009 D
V11 P010 N016 1.03
V12 N010 P009 1
D13 REF P011 D
D14 P012 REF D
V13 P012 VNEGx .3
V14 VPOSx P011 .3
D15 N013 P013 D
D16 P014 N013 D
V15 P014 VNEGx 0.6
V16 VPOSx P013 0.6
E4 Inverting_Out 0 N003 0 1
E5 noninverting_out 0 N012 0 1
Q1 Inv_Fdbk N002 RG- 0 PNP
Q2 Pos_Fdbk N015 RG+ 0 PNP
V1 VBIAS -Vs -10
I1 Pos_Fdbk VBIAS 9E-6
I2 Inv_Fdbk VBIAS 9E-6

C1 N003 Inv_Fdbk 3.8035e-12
C2 N012 Pos_Fdbk 3.8e-12
E8 N002 0 N005 0 1
E9 N015 0 N019 0 1
VOSI_Neg N004 IN- 25E-6
VOSI_Pos IN+ N017 24E-6
VOSO VOUT N011 300E-6
C3 RG- 0 .200e-12
C4 RG+ 0 .135e-12
I23 IN- 0 3E-12
I24 IN+ 0 3.2E-12
G1 0 IN+ N020 N021 .7e-9
R13 IN+ N020 10e9
R14 N020 IN- 10e9
R15 +Vs N021 10e9
R16 N021 -Vs 10e9
G2 0 IN- N020 N021 .7e-9
E10 VPOSx 0 +Vs 0 1
I3 +Vs -Vs 725E-6
G3 +Vs -Vs +Vs -Vs 1e-6
E11 VNEGx 0 -Vs 0 1

R17 VBIAS Inv_Fdbk 10e9
R18 Pos_Fdbk VBIAS 10e9
H3 N006 N004 V24 14
V24 N001 0 0
R19 N001 0 .0166
H4 N011 N009 V25 100
V25 N007 0 0
R20 N007 0 .0166
H5 N018 N017 V26 14
V26 N014 0 0
R21 N014 0 .0166
G4 0 N005 N006 N005 1E-3
G5 0 N019 N018 N019 1E-3
G6 0 N003 VBIAS Inv_Fdbk 1
G7 0 N012 VBIAS Pos_Fdbk 1
G8 0 N009 N013 N008 1
R10 N005 0 10e9
R7 N003 0 10E9
R11 N019 0 10E9
R8 N012 0 10E9
R9 N009 0 10E9
*C5 N008 N009 8e-12


H1 VPOSx N010 POLY(1) VOSO 0 0 8000
H2 N016 VNEGx POLY(1) VOSO 0 0 8000

* MODELS USED
*
.model D D
.model PNP PNP (BF=10E5 VAF=20000)
.ENDS AD8220

